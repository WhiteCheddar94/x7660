// ELEX 7660 Lab 4 
// Nicholas Scott AKA "White Cheddar"
// A01255181
// Feb. 6th, 2024
// Instructor: Sweet Bobby T

